// jtag_uart.v

// Generated using ACDS version 13.0sp1 232 at 2020.07.17.11:24:51

`timescale 1 ps / 1 ps
module jtag_uart (
		input  wire        clk_clk,                   //           clk.clk
		input  wire        reset_reset_n,             //         reset.reset_n
		input  wire        avbus_w8_r64_chipselect,   //  avbus_w8_r64.chipselect
		input  wire        avbus_w8_r64_address,      //              .address
		input  wire        avbus_w8_r64_read_n,       //              .read_n
		output wire [31:0] avbus_w8_r64_readdata,     //              .readdata
		input  wire        avbus_w8_r64_write_n,      //              .write_n
		input  wire [31:0] avbus_w8_r64_writedata,    //              .writedata
		output wire        avbus_w8_r64_waitrequest,  //              .waitrequest
		input  wire        avbus_w16_r32_chipselect,  // avbus_w16_r32.chipselect
		input  wire        avbus_w16_r32_address,     //              .address
		input  wire        avbus_w16_r32_read_n,      //              .read_n
		output wire [31:0] avbus_w16_r32_readdata,    //              .readdata
		input  wire        avbus_w16_r32_write_n,     //              .write_n
		input  wire [31:0] avbus_w16_r32_writedata,   //              .writedata
		output wire        avbus_w16_r32_waitrequest, //              .waitrequest
		input  wire        avbus_w32r16_chipselect,   //  avbus_w32r16.chipselect
		input  wire        avbus_w32r16_address,      //              .address
		input  wire        avbus_w32r16_read_n,       //              .read_n
		output wire [31:0] avbus_w32r16_readdata,     //              .readdata
		input  wire        avbus_w32r16_write_n,      //              .write_n
		input  wire [31:0] avbus_w32r16_writedata,    //              .writedata
		output wire        avbus_w32r16_waitrequest   //              .waitrequest
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [jtag_uart_w16_r32:rst_n, jtag_uart_w32_r8:rst_n, jtag_uart_w8_r64:rst_n]

	jtag_uart_jtag_uart_w16_r32 jtag_uart_w16_r32 (
		.clk            (clk_clk),                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset), //             reset.reset_n
		.av_chipselect  (avbus_w16_r32_chipselect),        // avalon_jtag_slave.chipselect
		.av_address     (avbus_w16_r32_address),           //                  .address
		.av_read_n      (avbus_w16_r32_read_n),            //                  .read_n
		.av_readdata    (avbus_w16_r32_readdata),          //                  .readdata
		.av_write_n     (avbus_w16_r32_write_n),           //                  .write_n
		.av_writedata   (avbus_w16_r32_writedata),         //                  .writedata
		.av_waitrequest (avbus_w16_r32_waitrequest),       //                  .waitrequest
		.av_irq         ()                                 //               irq.irq
	);

	jtag_uart_jtag_uart_w8_r64 jtag_uart_w8_r64 (
		.clk            (clk_clk),                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset), //             reset.reset_n
		.av_chipselect  (avbus_w8_r64_chipselect),         // avalon_jtag_slave.chipselect
		.av_address     (avbus_w8_r64_address),            //                  .address
		.av_read_n      (avbus_w8_r64_read_n),             //                  .read_n
		.av_readdata    (avbus_w8_r64_readdata),           //                  .readdata
		.av_write_n     (avbus_w8_r64_write_n),            //                  .write_n
		.av_writedata   (avbus_w8_r64_writedata),          //                  .writedata
		.av_waitrequest (avbus_w8_r64_waitrequest),        //                  .waitrequest
		.av_irq         ()                                 //               irq.irq
	);

	jtag_uart_jtag_uart_w32_r8 jtag_uart_w32_r8 (
		.clk            (clk_clk),                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset), //             reset.reset_n
		.av_chipselect  (avbus_w32r16_chipselect),         // avalon_jtag_slave.chipselect
		.av_address     (avbus_w32r16_address),            //                  .address
		.av_read_n      (avbus_w32r16_read_n),             //                  .read_n
		.av_readdata    (avbus_w32r16_readdata),           //                  .readdata
		.av_write_n     (avbus_w32r16_write_n),            //                  .write_n
		.av_writedata   (avbus_w32r16_writedata),          //                  .writedata
		.av_waitrequest (avbus_w32r16_waitrequest),        //                  .waitrequest
		.av_irq         ()                                 //               irq.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
