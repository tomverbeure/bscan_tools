// jtag_uart.v

// Generated using ACDS version 13.0sp1 232 at 2020.07.19.19:28:52

`timescale 1 ps / 1 ps
module jtag_uart (
		input  wire        clk_clk,           //   clk.clk
		input  wire        reset_reset_n,     // reset.reset_n
		input  wire        avbus_chipselect,  // avbus.chipselect
		input  wire        avbus_address,     //      .address
		input  wire        avbus_read_n,      //      .read_n
		output wire [31:0] avbus_readdata,    //      .readdata
		input  wire        avbus_write_n,     //      .write_n
		input  wire [31:0] avbus_writedata,   //      .writedata
		output wire        avbus_waitrequest  //      .waitrequest
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> jtag_uart_w8_r8:rst_n

	jtag_uart_jtag_uart_w8_r8 jtag_uart_w8_r8 (
		.clk            (clk_clk),                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset), //             reset.reset_n
		.av_chipselect  (avbus_chipselect),                // avalon_jtag_slave.chipselect
		.av_address     (avbus_address),                   //                  .address
		.av_read_n      (avbus_read_n),                    //                  .read_n
		.av_readdata    (avbus_readdata),                  //                  .readdata
		.av_write_n     (avbus_write_n),                   //                  .write_n
		.av_writedata   (avbus_writedata),                 //                  .writedata
		.av_waitrequest (avbus_waitrequest),               //                  .waitrequest
		.av_irq         ()                                 //               irq.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
